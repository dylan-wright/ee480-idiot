/*  
 *  EE480 - Assignment 2: The Making Of An IDIOT
 *  proccesor.v - top level module
 *  Version:
 *      03-02 : initial version
 *
 */

`define ALUadd 3'b000
`define ALUsub 3'b001
`define ALUxor 3'b010
`define ALUslt 3'b011
`define ALUor  3'b100
`define ALUand 3'b101
`define ALUsll 3'b110
`define ALUsrl 3'b111

module proccesor (
    input reset
    );

endmodule
