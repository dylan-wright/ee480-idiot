`include "signals.v"

module register_file(reg_out, reg_sel);
    input [5:0] reg_sel;
    output `WORD reg_out;

    reg registers[[[[[[[[[

endmodule
