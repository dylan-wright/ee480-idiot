module register_file(
