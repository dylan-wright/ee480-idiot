/*  
 *  EE480 - Assignment 2: The Making Of An IDIOT
 *  proccesor.v - top level module
 *  Version:
 *      03-02 : initial version
 *
 */

`include signals.v

module alu();
    input [WORD] X;
    input Y;
    
    output Z;

endmodule
