module dummy (
    input reset,
    output 
